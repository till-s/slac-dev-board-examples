library ieee;
use     ieee.std_logic_1164.all;
use     ieee.numeric_std.all;

use     work.ESCBasicTypesPkg.all;
use     work.Lan9254Pkg.all;
use     work.EEPROMConfigPkg.all;
use     work.EvrTxPDOPkg.all;

entity EEPROMConfiguratorTb is
end entity EEPROMConfiguratorTb;

architecture sim of EEPROMConfiguratorTb is

   constant SIZE_BYTES_C         : natural   := 2048;
   constant MAX_TXPDO_MAPS_C     : natural   := 16;

   signal clk                    : std_logic := '0';
   signal rst                    : std_logic := '1';

   signal sda                    : std_logic;
   signal scl                    : std_logic;
   signal scl_m_o                : std_logic;
   signal scl_m_t                : std_logic;
   signal sda_m_o                : std_logic;
   signal sda_m_t                : std_logic;
   signal scl_s_o                : std_logic := '1';
   signal sda_s_o                : std_logic := '1';

   signal run                    : boolean := true;

   signal ack                    : EEPROMConfigAckType := EEPROM_CONFIG_ACK_ASSERT_C;
   signal cfg                    : EEPROMConfigReqType;

   signal dbufMaps               : MemXferArray(MAX_TXPDO_MAPS_C - 1 downto 0);

   function toSlv(x : in Slv08Array) return std_logic_vector is
      variable v : std_logic_vector(8*x'length - 1 downto 0);
   begin
      for i in 0 to x'length - 1 loop
         v(8*i+7 downto 8*i) := x(x'low + i);
      end loop;
      return v;
   end function toSlv;

   constant EEPROM_INIT_0_C : Slv08Array(SIZE_BYTES_C - 1 downto 0) := (

      128    => x"51",
      129    => x"00",
      130    => std_logic_vector( to_unsigned( (160 - 128 - 4) / 2, 8 ) ),
      131    => x"00",
      132    => x"80",
      133    => x"10",
      134    => x"01",
      135    => x"00",

      160    => x"50",
      161    => x"00",
      162    => std_logic_vector( to_unsigned( (170 - 160 - 4) / 2, 8 ) ),
      163    => x"00",
      164    => x"00",
      165    => x"aa",
      166    => x"21",
      167    => x"43",

      170    => x"31", -- sync-manager
      171    => x"00",
      172    => std_logic_vector( to_unsigned( (256 - 170 - 2*4)/2, 8) ),
      173    => x"00",

      174 + 2*8 + 2 => x"04", -- SM2 length
      174 + 2*8 + 3 => x"00",

      174 + 3*8 + 2 => x"88", -- SM3 length
      174 + 3*8 + 3 => x"00",


      252    => x"01", -- category header
      253    => x"00", --
      254    => x"20", -- size (words)
      255    => x"00", --

      256    => x"56", -- mac addr
      257    => x"01",
      258    => x"02",
      259    => x"03",
      260    => x"04",
      261    => x"05",

      262    => x"0a", -- ip addr
      263    => x"0b",
      264    => x"0c",
      265    => x"0d",

      266    => x"40", -- udp port
      267    => x"50",

      268    => x"11", -- txPDO elements
      269    => x"00", -- ignored

      270    => x"04", -- txPDO mapping 0
      271    => x"20",
      272    => x"ef",
      273    => x"be",

      274    => x"00", -- txPDO mapping 1
      275    => x"01",
      276    => x"fe",
      277    => x"ca",
      others => x"FF"
   );

   constant EEPROM_INIT_1_C : Slv08Array(SIZE_BYTES_C - 1 downto 0) := (
      16#00000000# => x"91",
      16#00000001# => x"02",
      16#00000002# => x"01",
      16#00000003# => x"44",
      16#00000004# => x"00",
      16#00000005# => x"00",
      16#00000006# => x"00",
      16#00000007# => x"00",
      16#00000008# => x"00",
      16#00000009# => x"00",
      16#0000000a# => x"00",
      16#0000000b# => x"40",
      16#0000000c# => x"00",
      16#0000000d# => x"00",
      16#0000000e# => x"2b",
      16#0000000f# => x"00",
      16#00000010# => x"37",
      16#00000011# => x"13",
      16#00000012# => x"00",
      16#00000013# => x"00",
      16#00000014# => x"d2",
      16#00000015# => x"04",
      16#00000016# => x"00",
      16#00000017# => x"00",
      16#00000018# => x"00",
      16#00000019# => x"00",
      16#0000001a# => x"00",
      16#0000001b# => x"00",
      16#0000001c# => x"00",
      16#0000001d# => x"00",
      16#0000001e# => x"00",
      16#0000001f# => x"00",
      16#00000020# => x"00",
      16#00000021# => x"00",
      16#00000022# => x"00",
      16#00000023# => x"00",
      16#00000024# => x"00",
      16#00000025# => x"00",
      16#00000026# => x"00",
      16#00000027# => x"00",
      16#00000028# => x"00",
      16#00000029# => x"10",
      16#0000002a# => x"80",
      16#0000002b# => x"00",
      16#0000002c# => x"80",
      16#0000002d# => x"10",
      16#0000002e# => x"80",
      16#0000002f# => x"00",
      16#00000030# => x"00",
      16#00000031# => x"10",
      16#00000032# => x"30",
      16#00000033# => x"00",
      16#00000034# => x"80",
      16#00000035# => x"10",
      16#00000036# => x"30",
      16#00000037# => x"00",
      16#00000038# => x"22",
      16#00000039# => x"00",
      16#0000003a# => x"00",
      16#0000003b# => x"00",
      16#0000003c# => x"00",
      16#0000003d# => x"00",
      16#0000003e# => x"00",
      16#0000003f# => x"00",
      16#00000040# => x"00",
      16#00000041# => x"00",
      16#00000042# => x"00",
      16#00000043# => x"00",
      16#00000044# => x"00",
      16#00000045# => x"00",
      16#00000046# => x"00",
      16#00000047# => x"00",
      16#00000048# => x"00",
      16#00000049# => x"00",
      16#0000004a# => x"00",
      16#0000004b# => x"00",
      16#0000004c# => x"00",
      16#0000004d# => x"00",
      16#0000004e# => x"00",
      16#0000004f# => x"00",
      16#00000050# => x"00",
      16#00000051# => x"00",
      16#00000052# => x"00",
      16#00000053# => x"00",
      16#00000054# => x"00",
      16#00000055# => x"00",
      16#00000056# => x"00",
      16#00000057# => x"00",
      16#00000058# => x"00",
      16#00000059# => x"00",
      16#0000005a# => x"00",
      16#0000005b# => x"00",
      16#0000005c# => x"00",
      16#0000005d# => x"00",
      16#0000005e# => x"00",
      16#0000005f# => x"00",
      16#00000060# => x"00",
      16#00000061# => x"00",
      16#00000062# => x"00",
      16#00000063# => x"00",
      16#00000064# => x"00",
      16#00000065# => x"00",
      16#00000066# => x"00",
      16#00000067# => x"00",
      16#00000068# => x"00",
      16#00000069# => x"00",
      16#0000006a# => x"00",
      16#0000006b# => x"00",
      16#0000006c# => x"00",
      16#0000006d# => x"00",
      16#0000006e# => x"00",
      16#0000006f# => x"00",
      16#00000070# => x"00",
      16#00000071# => x"00",
      16#00000072# => x"00",
      16#00000073# => x"00",
      16#00000074# => x"00",
      16#00000075# => x"00",
      16#00000076# => x"00",
      16#00000077# => x"00",
      16#00000078# => x"00",
      16#00000079# => x"00",
      16#0000007a# => x"00",
      16#0000007b# => x"00",
      16#0000007c# => x"0f",
      16#0000007d# => x"00",
      16#0000007e# => x"01",
      16#0000007f# => x"00",
      16#00000080# => x"01",
      16#00000081# => x"00",
      16#00000082# => x"06",
      16#00000083# => x"00",
      16#00000084# => x"48",
      16#00000085# => x"02",
      16#00000086# => x"03",
      16#00000087# => x"04",
      16#00000088# => x"05",
      16#00000089# => x"66",
      16#0000008a# => x"00",
      16#0000008b# => x"00",
      16#0000008c# => x"00",
      16#0000008d# => x"00",
      16#0000008e# => x"00",
      16#0000008f# => x"00",
      16#00000090# => x"0a",
      16#00000091# => x"00",
      16#00000092# => x"1a",
      16#00000093# => x"00",
      16#00000094# => x"07",
      16#00000095# => x"0b",
      16#00000096# => x"6c",
      16#00000097# => x"61",
      16#00000098# => x"6e",
      16#00000099# => x"39",
      16#0000009a# => x"32",
      16#0000009b# => x"35",
      16#0000009c# => x"32",
      16#0000009d# => x"5f",
      16#0000009e# => x"73",
      16#0000009f# => x"70",
      16#000000a0# => x"69",
      16#000000a1# => x"07",
      16#000000a2# => x"6c",
      16#000000a3# => x"61",
      16#000000a4# => x"6e",
      16#000000a5# => x"39",
      16#000000a6# => x"32",
      16#000000a7# => x"35",
      16#000000a8# => x"32",
      16#000000a9# => x"04",
      16#000000aa# => x"4c",
      16#000000ab# => x"45",
      16#000000ac# => x"44",
      16#000000ad# => x"73",
      16#000000ae# => x"04",
      16#000000af# => x"4c",
      16#000000b0# => x"45",
      16#000000b1# => x"44",
      16#000000b2# => x"30",
      16#000000b3# => x"04",
      16#000000b4# => x"4c",
      16#000000b5# => x"45",
      16#000000b6# => x"44",
      16#000000b7# => x"31",
      16#000000b8# => x"07",
      16#000000b9# => x"42",
      16#000000ba# => x"75",
      16#000000bb# => x"74",
      16#000000bc# => x"74",
      16#000000bd# => x"6f",
      16#000000be# => x"6e",
      16#000000bf# => x"73",
      16#000000c0# => x"07",
      16#000000c1# => x"42",
      16#000000c2# => x"75",
      16#000000c3# => x"74",
      16#000000c4# => x"74",
      16#000000c5# => x"6f",
      16#000000c6# => x"6e",
      16#000000c7# => x"31",
      16#000000c8# => x"1e",
      16#000000c9# => x"00",
      16#000000ca# => x"10",
      16#000000cb# => x"00",
      16#000000cc# => x"01",
      16#000000cd# => x"00",
      16#000000ce# => x"00",
      16#000000cf# => x"02",
      16#000000d0# => x"00",
      16#000000d1# => x"00",
      16#000000d2# => x"00",
      16#000000d3# => x"01",
      16#000000d4# => x"00",
      16#000000d5# => x"00",
      16#000000d6# => x"00",
      16#000000d7# => x"00",
      16#000000d8# => x"00",
      16#000000d9# => x"00",
      16#000000da# => x"01",
      16#000000db# => x"00",
      16#000000dc# => x"11",
      16#000000dd# => x"00",
      16#000000de# => x"00",
      16#000000df# => x"00",
      16#000000e0# => x"00",
      16#000000e1# => x"00",
      16#000000e2# => x"00",
      16#000000e3# => x"00",
      16#000000e4# => x"00",
      16#000000e5# => x"00",
      16#000000e6# => x"00",
      16#000000e7# => x"00",
      16#000000e8# => x"00",
      16#000000e9# => x"00",
      16#000000ea# => x"00",
      16#000000eb# => x"00",
      16#000000ec# => x"28",
      16#000000ed# => x"00",
      16#000000ee# => x"01",
      16#000000ef# => x"00",
      16#000000f0# => x"01",
      16#000000f1# => x"02",
      16#000000f2# => x"29",
      16#000000f3# => x"00",
      16#000000f4# => x"10",
      16#000000f5# => x"00",
      16#000000f6# => x"00",
      16#000000f7# => x"10",
      16#000000f8# => x"30",
      16#000000f9# => x"00",
      16#000000fa# => x"26",
      16#000000fb# => x"00",
      16#000000fc# => x"01",
      16#000000fd# => x"01",
      16#000000fe# => x"80",
      16#000000ff# => x"10",
      16#00000100# => x"30",
      16#00000101# => x"00",
      16#00000102# => x"22",
      16#00000103# => x"00",
      16#00000104# => x"01",
      16#00000105# => x"02",
      16#00000106# => x"00",
      16#00000107# => x"11",
      16#00000108# => x"03",
      16#00000109# => x"00",
      16#0000010a# => x"24",
      16#0000010b# => x"00",
      16#0000010c# => x"01",
      16#0000010d# => x"03",
      16#0000010e# => x"80",
      16#0000010f# => x"11",
      16#00000110# => x"04",
      16#00000111# => x"00",
      16#00000112# => x"20",
      16#00000113# => x"00",
      16#00000114# => x"01",
      16#00000115# => x"04",
      16#00000116# => x"32",
      16#00000117# => x"00",
      16#00000118# => x"08",
      16#00000119# => x"00",
      16#0000011a# => x"00",
      16#0000011b# => x"1a",
      16#0000011c# => x"01",
      16#0000011d# => x"03",
      16#0000011e# => x"00",
      16#0000011f# => x"06",
      16#00000120# => x"00",
      16#00000121# => x"00",
      16#00000122# => x"00",
      16#00000123# => x"60",
      16#00000124# => x"01",
      16#00000125# => x"07",
      16#00000126# => x"01",
      16#00000127# => x"20",
      16#00000128# => x"00",
      16#00000129# => x"00",
      16#0000012a# => x"33",
      16#0000012b# => x"00",
      16#0000012c# => x"0c",
      16#0000012d# => x"00",
      16#0000012e# => x"00",
      16#0000012f# => x"16",
      16#00000130# => x"02",
      16#00000131# => x"02",
      16#00000132# => x"00",
      16#00000133# => x"03",
      16#00000134# => x"00",
      16#00000135# => x"00",
      16#00000136# => x"00",
      16#00000137# => x"70",
      16#00000138# => x"01",
      16#00000139# => x"04",
      16#0000013a# => x"01",
      16#0000013b# => x"08",
      16#0000013c# => x"00",
      16#0000013d# => x"00",
      16#0000013e# => x"00",
      16#0000013f# => x"70",
      16#00000140# => x"02",
      16#00000141# => x"05",
      16#00000142# => x"01",
      16#00000143# => x"08",
      16#00000144# => x"00",
      16#00000145# => x"00",
      16#00000146# => x"ff",
      16#00000147# => x"ff",
      others    => (others => '1')
   );

   constant EEPROM_INIT_2_C : Slv08Array(SIZE_BYTES_C - 1 downto 0) := (
   0 => x"91",
   1 => x"02",
   2 => x"01",
   3 => x"44",
   4 => x"00",
   5 => x"00",
   6 => x"00",
   7 => x"00",
   8 => x"00",
   9 => x"00",
   10 => x"00",
   11 => x"40",
   12 => x"00",
   13 => x"00",
   14 => x"2b",
   15 => x"00",
   16 => x"49",
   17 => x"53",
   18 => x"50",
   19 => x"00",
   20 => x"01",
   21 => x"00",
   22 => x"00",
   23 => x"00",
   24 => x"01",
   25 => x"00",
   26 => x"00",
   27 => x"00",
   28 => x"00",
   29 => x"00",
   30 => x"00",
   31 => x"00",
   32 => x"00",
   33 => x"00",
   34 => x"00",
   35 => x"00",
   36 => x"00",
   37 => x"00",
   38 => x"00",
   39 => x"00",
   40 => x"00",
   41 => x"00",
   42 => x"00",
   43 => x"00",
   44 => x"00",
   45 => x"00",
   46 => x"00",
   47 => x"00",
   48 => x"00",
   49 => x"10",
   50 => x"30",
   51 => x"00",
   52 => x"80",
   53 => x"10",
   54 => x"30",
   55 => x"00",
   56 => x"02",
   57 => x"00",
   58 => x"00",
   59 => x"00",
   60 => x"00",
   61 => x"00",
   62 => x"00",
   63 => x"00",
   64 => x"00",
   65 => x"00",
   66 => x"00",
   67 => x"00",
   68 => x"00",
   69 => x"00",
   70 => x"00",
   71 => x"00",
   72 => x"00",
   73 => x"00",
   74 => x"00",
   75 => x"00",
   76 => x"00",
   77 => x"00",
   78 => x"00",
   79 => x"00",
   80 => x"00",
   81 => x"00",
   82 => x"00",
   83 => x"00",
   84 => x"00",
   85 => x"00",
   86 => x"00",
   87 => x"00",
   88 => x"00",
   89 => x"00",
   90 => x"00",
   91 => x"00",
   92 => x"00",
   93 => x"00",
   94 => x"00",
   95 => x"00",
   96 => x"00",
   97 => x"00",
   98 => x"00",
   99 => x"00",
   100 => x"00",
   101 => x"00",
   102 => x"00",
   103 => x"00",
   104 => x"00",
   105 => x"00",
   106 => x"00",
   107 => x"00",
   108 => x"00",
   109 => x"00",
   110 => x"00",
   111 => x"00",
   112 => x"00",
   113 => x"00",
   114 => x"00",
   115 => x"00",
   116 => x"00",
   117 => x"00",
   118 => x"00",
   119 => x"00",
   120 => x"00",
   121 => x"00",
   122 => x"00",
   123 => x"00",
   124 => x"0f",
   125 => x"00",
   126 => x"01",
   127 => x"00",
   128 => x"01",
   129 => x"00",
   130 => x"07",
   131 => x"00",
   132 => x"48",
   133 => x"01",
   134 => x"02",
   135 => x"03",
   136 => x"04",
   137 => x"05",
   138 => x"0a",
   139 => x"0a",
   140 => x"0a",
   141 => x"0b",
   142 => x"ff",
   143 => x"ff",
   144 => x"3f",
   145 => x"00",
   146 => x"0a",
   147 => x"00",
   148 => x"7d",
   149 => x"00",
   150 => x"14",
   151 => x"07",
   152 => x"4c",
   153 => x"61",
   154 => x"6e",
   155 => x"39",
   156 => x"32",
   157 => x"35",
   158 => x"34",
   159 => x"05",
   160 => x"45",
   161 => x"63",
   162 => x"45",
   163 => x"56",
   164 => x"52",
   165 => x"06",
   166 => x"4c",
   167 => x"45",
   168 => x"44",
   169 => x"5b",
   170 => x"30",
   171 => x"5d",
   172 => x"06",
   173 => x"4c",
   174 => x"45",
   175 => x"44",
   176 => x"5b",
   177 => x"31",
   178 => x"5d",
   179 => x"06",
   180 => x"4c",
   181 => x"45",
   182 => x"44",
   183 => x"5b",
   184 => x"32",
   185 => x"5d",
   186 => x"13",
   187 => x"45",
   188 => x"43",
   189 => x"41",
   190 => x"54",
   191 => x"20",
   192 => x"45",
   193 => x"56",
   194 => x"52",
   195 => x"20",
   196 => x"44",
   197 => x"61",
   198 => x"74",
   199 => x"61",
   200 => x"62",
   201 => x"75",
   202 => x"66",
   203 => x"66",
   204 => x"65",
   205 => x"72",
   206 => x"0b",
   207 => x"54",
   208 => x"69",
   209 => x"6d",
   210 => x"65",
   211 => x"73",
   212 => x"74",
   213 => x"61",
   214 => x"6d",
   215 => x"70",
   216 => x"48",
   217 => x"69",
   218 => x"0b",
   219 => x"54",
   220 => x"69",
   221 => x"6d",
   222 => x"65",
   223 => x"73",
   224 => x"74",
   225 => x"61",
   226 => x"6d",
   227 => x"70",
   228 => x"4c",
   229 => x"6f",
   230 => x"09",
   231 => x"45",
   232 => x"76",
   233 => x"65",
   234 => x"6e",
   235 => x"74",
   236 => x"73",
   237 => x"5b",
   238 => x"30",
   239 => x"5d",
   240 => x"09",
   241 => x"45",
   242 => x"76",
   243 => x"65",
   244 => x"6e",
   245 => x"74",
   246 => x"73",
   247 => x"5b",
   248 => x"31",
   249 => x"5d",
   250 => x"09",
   251 => x"45",
   252 => x"76",
   253 => x"65",
   254 => x"6e",
   255 => x"74",
   256 => x"73",
   257 => x"5b",
   258 => x"32",
   259 => x"5d",
   260 => x"09",
   261 => x"45",
   262 => x"76",
   263 => x"65",
   264 => x"6e",
   265 => x"74",
   266 => x"73",
   267 => x"5b",
   268 => x"33",
   269 => x"5d",
   270 => x"09",
   271 => x"45",
   272 => x"76",
   273 => x"65",
   274 => x"6e",
   275 => x"74",
   276 => x"73",
   277 => x"5b",
   278 => x"34",
   279 => x"5d",
   280 => x"09",
   281 => x"45",
   282 => x"76",
   283 => x"65",
   284 => x"6e",
   285 => x"74",
   286 => x"73",
   287 => x"5b",
   288 => x"35",
   289 => x"5d",
   290 => x"09",
   291 => x"45",
   292 => x"76",
   293 => x"65",
   294 => x"6e",
   295 => x"74",
   296 => x"73",
   297 => x"5b",
   298 => x"36",
   299 => x"5d",
   300 => x"09",
   301 => x"45",
   302 => x"76",
   303 => x"65",
   304 => x"6e",
   305 => x"74",
   306 => x"73",
   307 => x"5b",
   308 => x"37",
   309 => x"5d",
   310 => x"15",
   311 => x"54",
   312 => x"69",
   313 => x"6d",
   314 => x"65",
   315 => x"73",
   316 => x"74",
   317 => x"61",
   318 => x"6d",
   319 => x"70",
   320 => x"4c",
   321 => x"61",
   322 => x"74",
   323 => x"63",
   324 => x"68",
   325 => x"30",
   326 => x"52",
   327 => x"69",
   328 => x"73",
   329 => x"69",
   330 => x"6e",
   331 => x"67",
   332 => x"16",
   333 => x"54",
   334 => x"69",
   335 => x"6d",
   336 => x"65",
   337 => x"73",
   338 => x"74",
   339 => x"61",
   340 => x"6d",
   341 => x"70",
   342 => x"4c",
   343 => x"61",
   344 => x"74",
   345 => x"63",
   346 => x"68",
   347 => x"30",
   348 => x"46",
   349 => x"61",
   350 => x"6c",
   351 => x"6c",
   352 => x"69",
   353 => x"6e",
   354 => x"67",
   355 => x"15",
   356 => x"54",
   357 => x"69",
   358 => x"6d",
   359 => x"65",
   360 => x"73",
   361 => x"74",
   362 => x"61",
   363 => x"6d",
   364 => x"70",
   365 => x"4c",
   366 => x"61",
   367 => x"74",
   368 => x"63",
   369 => x"68",
   370 => x"31",
   371 => x"52",
   372 => x"69",
   373 => x"73",
   374 => x"69",
   375 => x"6e",
   376 => x"67",
   377 => x"16",
   378 => x"54",
   379 => x"69",
   380 => x"6d",
   381 => x"65",
   382 => x"73",
   383 => x"74",
   384 => x"61",
   385 => x"6d",
   386 => x"70",
   387 => x"4c",
   388 => x"61",
   389 => x"74",
   390 => x"63",
   391 => x"68",
   392 => x"31",
   393 => x"46",
   394 => x"61",
   395 => x"6c",
   396 => x"6c",
   397 => x"69",
   398 => x"6e",
   399 => x"67",
   400 => x"1e",
   401 => x"00",
   402 => x"10",
   403 => x"00",
   404 => x"01",
   405 => x"00",
   406 => x"00",
   407 => x"02",
   408 => x"00",
   409 => x"00",
   410 => x"00",
   411 => x"01",
   412 => x"00",
   413 => x"00",
   414 => x"00",
   415 => x"00",
   416 => x"00",
   417 => x"00",
   418 => x"01",
   419 => x"00",
   420 => x"11",
   421 => x"00",
   422 => x"00",
   423 => x"00",
   424 => x"00",
   425 => x"00",
   426 => x"00",
   427 => x"00",
   428 => x"00",
   429 => x"00",
   430 => x"00",
   431 => x"00",
   432 => x"00",
   433 => x"00",
   434 => x"00",
   435 => x"00",
   436 => x"28",
   437 => x"00",
   438 => x"02",
   439 => x"00",
   440 => x"02",
   441 => x"01",
   442 => x"00",
   443 => x"00",
   444 => x"29",
   445 => x"00",
   446 => x"10",
   447 => x"00",
   448 => x"00",
   449 => x"10",
   450 => x"30",
   451 => x"00",
   452 => x"26",
   453 => x"00",
   454 => x"01",
   455 => x"01",
   456 => x"80",
   457 => x"10",
   458 => x"30",
   459 => x"00",
   460 => x"22",
   461 => x"00",
   462 => x"01",
   463 => x"02",
   464 => x"00",
   465 => x"11",
   466 => x"03",
   467 => x"00",
   468 => x"24",
   469 => x"00",
   470 => x"01",
   471 => x"03",
   472 => x"80",
   473 => x"11",
   474 => x"48",
   475 => x"00",
   476 => x"20",
   477 => x"00",
   478 => x"01",
   479 => x"04",
   480 => x"32",
   481 => x"00",
   482 => x"3c",
   483 => x"00",
   484 => x"00",
   485 => x"1a",
   486 => x"0e",
   487 => x"03",
   488 => x"00",
   489 => x"06",
   490 => x"00",
   491 => x"00",
   492 => x"00",
   493 => x"50",
   494 => x"01",
   495 => x"07",
   496 => x"07",
   497 => x"20",
   498 => x"00",
   499 => x"00",
   500 => x"01",
   501 => x"50",
   502 => x"01",
   503 => x"08",
   504 => x"07",
   505 => x"20",
   506 => x"00",
   507 => x"00",
   508 => x"02",
   509 => x"50",
   510 => x"01",
   511 => x"09",
   512 => x"07",
   513 => x"20",
   514 => x"00",
   515 => x"00",
   516 => x"02",
   517 => x"50",
   518 => x"02",
   519 => x"0a",
   520 => x"07",
   521 => x"20",
   522 => x"00",
   523 => x"00",
   524 => x"02",
   525 => x"50",
   526 => x"03",
   527 => x"0b",
   528 => x"07",
   529 => x"20",
   530 => x"00",
   531 => x"00",
   532 => x"02",
   533 => x"50",
   534 => x"04",
   535 => x"0c",
   536 => x"07",
   537 => x"20",
   538 => x"00",
   539 => x"00",
   540 => x"02",
   541 => x"50",
   542 => x"05",
   543 => x"0d",
   544 => x"07",
   545 => x"20",
   546 => x"00",
   547 => x"00",
   548 => x"02",
   549 => x"50",
   550 => x"06",
   551 => x"0e",
   552 => x"07",
   553 => x"20",
   554 => x"00",
   555 => x"00",
   556 => x"02",
   557 => x"50",
   558 => x"07",
   559 => x"0f",
   560 => x"07",
   561 => x"20",
   562 => x"00",
   563 => x"00",
   564 => x"02",
   565 => x"50",
   566 => x"08",
   567 => x"10",
   568 => x"07",
   569 => x"20",
   570 => x"00",
   571 => x"00",
   572 => x"03",
   573 => x"50",
   574 => x"01",
   575 => x"11",
   576 => x"1b",
   577 => x"40",
   578 => x"00",
   579 => x"00",
   580 => x"04",
   581 => x"50",
   582 => x"01",
   583 => x"12",
   584 => x"1b",
   585 => x"40",
   586 => x"00",
   587 => x"00",
   588 => x"05",
   589 => x"50",
   590 => x"01",
   591 => x"13",
   592 => x"1b",
   593 => x"40",
   594 => x"00",
   595 => x"00",
   596 => x"06",
   597 => x"50",
   598 => x"01",
   599 => x"14",
   600 => x"1b",
   601 => x"40",
   602 => x"00",
   603 => x"00",
   604 => x"33",
   605 => x"00",
   606 => x"10",
   607 => x"00",
   608 => x"00",
   609 => x"00",
   610 => x"03",
   611 => x"02",
   612 => x"00",
   613 => x"00",
   614 => x"00",
   615 => x"00",
   616 => x"00",
   617 => x"20",
   618 => x"01",
   619 => x"03",
   620 => x"05",
   621 => x"08",
   622 => x"00",
   623 => x"00",
   624 => x"00",
   625 => x"20",
   626 => x"02",
   627 => x"04",
   628 => x"05",
   629 => x"08",
   630 => x"00",
   631 => x"00",
   632 => x"00",
   633 => x"20",
   634 => x"03",
   635 => x"05",
   636 => x"05",
   637 => x"08",
   638 => x"00",
   639 => x"00",
   640 => x"ff",
   641 => x"ff",
   others => x"ff"
   );

   constant EEPROM_INIT_C : Slv08Array := EEPROM_INIT_2_C;

begin

   sda <= (sda_m_t or sda_m_o) and sda_s_o;
   scl <= (scl_m_t or scl_m_o) and scl_s_o;

   P_CLK : process is
   begin
      if ( run ) then
         wait for 1.25 us;
         clk <= not clk;
      else
         wait;
      end if;
   end process P_CLK;

   P_DRV : process is
   begin
      wait until rising_edge( clk );
      wait until rising_edge( clk );
      wait until rising_edge( clk );
      rst <= '0';
      wait until rising_edge( clk );
      wait;
   end process P_DRV;

   P_DON : process (clk) is
   begin
      if ( rising_edge( clk ) ) then
         if ( cfg.net.macAddrVld = '1' ) then
            report "MAC: " & toString( cfg.net.macAddr );
         end if;
         if ( cfg.net.ip4AddrVld = '1' ) then
            report "IP4: " & toString( cfg.net.ip4Addr );
         end if;
         if ( cfg.net.udpPortVld = '1' ) then
            report "UDP: " & toString( cfg.net.udpPort );
         end if;
         if ( cfg.esc.valid = '1' ) then
            report "NMAPS:   " & integer'image( cfg.txPDO.numMaps );
            report "SM2 LEN: " & toString( cfg.esc.sm2Len );
            report "SM3 LEN: " & toString( cfg.esc.sm3Len );
            for j in 0 to cfg.txPDO.numMaps - 1 loop
               report "MAP " & integer'image(j) & " : off " & toString( dbufMaps(j).off )
                                                & " : swp " & toString( dbufMaps(j).swp )
                                                & " : num " & toString( dbufMaps(j).num );
            end loop;
            report "DONE";
            run <= false;
         end if;
      end if;
   end process P_DON;

   U_EEP : entity work.I2CEEPROM
      generic map (
         SIZE_BYTES_G  => SIZE_BYTES_C,
         EEPROM_INIT_G => toSlv( EEPROM_INIT_C )
      )
      port map (
         clk       => clk,
         rst       => rst,

         sclSync   => scl,
         sdaSync   => sda,
         sdaOut    => sda_s_o
      );

   -- ClockFrequency_g must be >= 12*I2cFrequency_g
   -- otherwise spurious arbitration-lost will be detected
   -- (probably due to synchronizer delays)
   U_DUT : entity work.EEPROMConfigurator
      generic map (
         CLOCK_FREQ_G               => 5.0e5,
         I2C_FREQ_G                 => 4.0e4,
         EEPROM_OFFSET_G            => 0, --128,
         EEPROM_SIZE_G              => (8*SIZE_BYTES_C),
         MAX_TXPDO_MAPS_G           => MAX_TXPDO_MAPS_C,
         I2C_ADDR_G                 => "1010101"
      )
      port map (
         clk             => clk,
         rst             => rst,

         dbufMaps        => dbufMaps,
         configReq       => cfg,
         configAck       => ack,

         i2cSclInp       => scl,
         i2cSclOut       => scl_m_o,
         i2cSclHiZ       => scl_m_t,

         i2cSdaInp       => sda,
         i2cSdaOut       => sda_m_o,
         i2cSdaHiZ       => sda_m_t
      );
end architecture sim;

